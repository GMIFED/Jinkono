* On-die Decoupling circuit for V00H (VDDQ to VSSQ)
* Includes VDDQ-VSSQ decoupling for an individual signal such as DQ0-15, DQS, DQS#, or DM.
* This subcircuit should be added across the IBIS DQ, DM or DQS model's [Pullup Reference] and [Pulldown Reference]
* nodes as in the following Spice example:

******************************************************************************************************
*x_decouple vddq_die vssq_die v00h_ondie_decoupling_perdq

*b_dq1 vddq_die vssq_die PAD_DQ1 IN_DQ1 ENOUT RCVR_OUT_DQ1 vddq_die vssq_die 
*+ file='v00h_v5p0.ibs' model='DQ_34_2133' typ=typ power=off buffer=3 interpol=1 ramp_fwf=2 ramp_rwf=2
*+ rm_tail_rwf=default rm_tail_fwf=default
*+ rm_dly_rwf=default rm_dly_fwf=default
******************************************************************************************************


.subckt v00h_ondie_decoupling_perdq vddq_die vssq_die
x1 vddq_die vssq_die v00h_cfat_perdq



**********************************************************
** STATE-SPACE REALIZATION               
** IN SPICE LANGUAGE
** This file is automatically generated  
**********************************************************
** Created: 11-Aug-2015 by IdEM R2012 (8.0.6)
**********************************************************


**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt v00h_cfat_perdq
+  a_1 b_1 
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+001
GC_1_1 b_1 NI_1 NS_1 0 4.1865810284169809e-002
GC_1_2 b_1 NI_1 NS_2 0 2.2034190242812843e-003
GC_1_3 b_1 NI_1 NS_3 0 3.5300911213663888e-005
GC_1_4 b_1 NI_1 NS_4 0 1.1612512586435584e-005
GC_1_5 b_1 NI_1 NS_5 0 4.4163414864942093e-006
GC_1_6 b_1 NI_1 NS_6 0 2.0990549175006187e-004
GD_1_1 b_1 NI_1 NA_1 0 -2.8091649809949204e-001
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+000
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-002
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-013
RS_1 NS_1 0 3.9404233733066056e+000
GS_1_1 0 NS_1 NA_1 0 1.5673186053703178e-001
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-013
RS_2 NS_2 0 2.4563024341334931e+001
GS_2_1 0 NS_2 NA_1 0 1.5673186053703178e-001
*
* Real pole n. 3
CS_3 NS_3 0 9.9999999999999998e-013
RS_3 NS_3 0 3.8163796078901913e+002
GS_3_1 0 NS_3 NA_1 0 1.5673186053703178e-001
*
* Real pole n. 4
CS_4 NS_4 0 9.9999999999999998e-013
RS_4 NS_4 0 2.4441320188898972e+003
GS_4_1 0 NS_4 NA_1 0 1.5673186053703178e-001
*
* Real pole n. 5
CS_5 NS_5 0 9.9999999999999998e-013
RS_5 NS_5 0 3.3816169566555436e+004
GS_5_1 0 NS_5 NA_1 0 1.5673186053703178e-001
*
* Real pole n. 6
CS_6 NS_6 0 9.9999999999999998e-013
RS_6 NS_6 0 1.5179020843263068e+004
GS_6_1 0 NS_6 NA_1 0 1.5673186053703178e-001
*
******************************


.ends
*******************
* End of subcircuit
*******************
.ends
