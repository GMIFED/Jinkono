* On-die Decoupling circuit for V00H (VDDQ to VSSQ)
* Includes VDDQ-VSSQ decoupling for all signals (full die) including DDQ0-15, DQS, DQS#, or DM.
* This subcircuit should be added across the IBIS DQ and DQS models' [Pullup Reference] and [Pulldown Reference]
* nodes as in the following Spice example:

******************************************************************************************************
*x_decouple vddq_die vssq_die v00h_ondie_decoupling_all

*b_dq1 vddq_die vssq_die PAD_DQ1 IN_DQ1 ENOUT RCVR_OUT_DQ1 vddq_die vssq_die 
*+ file='v00h_v5p0.ibs' model='DQ_34_2133' typ=typ power=off buffer=3 interpol=1 ramp_fwf=2 ramp_rwf=2
*+ rm_tail_rwf=default rm_tail_fwf=default
*+ rm_dly_rwf=default rm_dly_fwf=default
******************************************************************************************************


.subckt v00h_ondie_decoupling_all vddq_die vssq_die
x1 vddq_die vssq_die v00h_cfat_all




**********************************************************
** STATE-SPACE REALIZATION               
** IN SPICE LANGUAGE
** This file is automatically generated  
**********************************************************
** Created: 11-Aug-2015 by IdEM R2012 (8.0.6)
**********************************************************


**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt v00h_cfat_all
+  a_1 b_1 
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+001
GC_1_1 b_1 NI_1 NS_1 0 2.5021483574124283e-003
GC_1_2 b_1 NI_1 NS_2 0 1.1049788915004628e-005
GC_1_3 b_1 NI_1 NS_3 0 4.4727021762869755e-007
GC_1_4 b_1 NI_1 NS_4 0 1.7339302549033419e-004
GD_1_1 b_1 NI_1 NA_1 0 -2.8170916819588471e-001
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+000
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-002
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-013
RS_1 NS_1 0 3.5619855263442162e+001
GS_1_1 0 NS_1 NA_1 0 9.5001155183608230e-003
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-013
RS_2 NS_2 0 1.0039094727016194e+005
GS_2_1 0 NS_2 NA_1 0 9.5001155183608230e-003
*
* Real pole n. 3
CS_3 NS_3 0 9.9999999999999998e-013
RS_3 NS_3 0 1.4354444876078407e+006
GS_3_1 0 NS_3 NA_1 0 9.5001155183608230e-003
*
* Real pole n. 4
CS_4 NS_4 0 9.9999999999999998e-013
RS_4 NS_4 0 3.3200946041646646e+005
GS_4_1 0 NS_4 NA_1 0 9.5001155183608230e-003
*
******************************


.ends
*******************
* End of subcircuit
*******************
.ends
